module network

#include <enet.h>

