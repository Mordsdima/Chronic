module engine

pub struct Context {

}