module main

import veb

pub fn (mut app App) profile_asset(mut ctx Context) veb.Result {
	return ctx.text('TODO')
}
