module types

pub struct Rect {
pub mut:
	x int
	y int
	w int
	h int
}