module network

