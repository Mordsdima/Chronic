module types

@[heap]
pub struct Context {
pub mut:
	r Renderer
}