module main

import network

fn main() {
	//network.init()
	println('Hello World!')
	
}
