module types

pub struct Rect {
pub mut:
	x f32
	y f32
	w f32
	h f32
}
