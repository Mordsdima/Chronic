module screens